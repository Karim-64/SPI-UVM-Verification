package SPI_wrapper_driver_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
import SPI_wrapper_config_pkg::*;
import SPI_wrapper_seq_item_pkg::*;
    class SPI_wrapper_driver extends uvm_driver #(SPI_wrapper_seq_item);
        `uvm_component_utils(SPI_wrapper_driver)
        virtual SPI_wrapper_if wrapper_vif;
        SPI_wrapper_seq_item stim_seq_item;

        function new(string name, uvm_component parent);
            super.new(name, parent);    
        endfunction

        task run_phase(uvm_phase phase);
            super.run_phase(phase);
            forever begin             
                stim_seq_item = SPI_wrapper_seq_item::type_id::create("stim_seq_item");
                seq_item_port.get_next_item(stim_seq_item);
                wrapper_vif.MOSI = stim_seq_item.MOSI;
                wrapper_vif.SS_n     = stim_seq_item.SS_n;
                wrapper_vif.rst_n = stim_seq_item.rst_n;
                @(negedge wrapper_vif.clk);
                seq_item_port.item_done();
            end
        endtask;
    endclass
endpackage