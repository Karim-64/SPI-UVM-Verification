package spi_slave_shared_pkg;
    parameter IDLE      = 3'b000;
    parameter WRITE     = 3'b001;
    parameter CHK_CMD   = 3'b010;
    parameter READ_ADD  = 3'b011;
    parameter READ_DATA = 3'b100;
endpackage